`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// Engineer: Dennis Hardy
// Module: MUL
//
//////////////////////////////////////////////////////////////////////////////////

module MUL #(parameter DATAWIDTH = 8) (a, b, prod);
   input [DATAWIDTH-1:0] a, b;

   output reg [2*DATAWIDTH-1:0] prod;

   always @ (a, b) begin
      prod <= a*b;
   end

endmodule // MUL
